

	`define SST_ON	//save state
	`define GGC_ON	//cheats engine
	`define SND_ON	//expansion sound if any exists
