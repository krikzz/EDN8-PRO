

module top
(cpu_dat, cpu_addr, cpu_ce, cpu_rw, cpu_m2, cpu_irq,
cpu_dir, cpu_ex,
spi_miso, spi_mosi, spi_clk, spi_ss,
ice_ss, ice_sck, ice_sdi, ice_sdo,
boot0, mcu_rst, 
clk, boot_on, gpio
);

	inout [7:0]cpu_dat;
	input [14:0]cpu_addr;
	input cpu_ce, cpu_rw, cpu_m2, cpu_irq;
	output cpu_dir, cpu_ex;

	
	output spi_miso;
	input spi_mosi, spi_clk, spi_ss;
	
	input ice_ss, ice_sck, ice_sdi;
	output ice_sdo;
	
	output boot0, mcu_rst;
	
	input clk, boot_on;
	output [3:0]gpio;
	
	
	assign cpu_dat[7:0] = 8'hzz;
	assign cpu_dir = boot_on ? 1 : 1'bz;
	assign cpu_ex =  boot_on ? !rom_oe : 1'bz;
	

	assign boot0 = 1'bz;
	assign mcu_rst = 1'bz;

	assign spi_miso = 1'bz;
	assign ice_sdo = 1'bz;
	
	assign gpio[3:0] = 4'bzzzz;
	
	assign cpu_dat[7:0] = rom_oe ? rom_dat[7:0] : 8'hzz;
	
	wire rom_oe = boot_on & cpu_rw & cpu_m2 & !cpu_ce;
	
	wire [7:0]rom_dat;
	
	boot1 rom_inst(clk, cpu_addr[9:0], rom_dat);
	
endmodule


module boot1(
	input clk,
	input [9:0]addr_rd_in,
	output [7:0]data_out
);

	

	defparam ram0.INIT_0 = 256'h20203030312E20766465636F6F74426F202020204E3865206976447265724576;
	defparam ram0.INIT_1 = 256'h6979736B6F7675626F6C20476F724967202049545A204B5A5249204B31393230;
	defparam ram0.INIT_2 = 256'h008DFBA920102C020220042C4C00D0F704E89D0055FC20BD8E00A200FF9A78A2;
	defparam ram0.INIT_3 = 256'h4908FF40FAADCAD00720208D0CA220A98D06A90006203F8D20A98D01A90A0020;
	defparam ram0.INIT_4 = 256'h06203F8DFBA920102C020220E82CA0D0F0C98A29D0EFC9012901F6AA40D0CDFF;
	defparam ram0.INIT_5 = 256'h0000000000000000000000004000FCFFFA6CCAD00720208D06A220A98D06A900;
	defparam ram0.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram0.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

	defparam ram1.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam ram1.INIT_F = 256'hB2FC40FCB2FC0000000000000000000000000000000000000000000000000000;

	wire [9:0]addr_rd = {addr_rd_in[9:1], !addr_rd_in[0]};
	assign data_out[7:0] = data_out_x[addr_rd[9]];
	wire [7:0]data_out_x[2];

	
	SB_RAM512x8NRNW ram0(
		.RDATA(data_out_x[0][7:0]),
		.RADDR(addr_rd[8:0]),
		.RCLKN(clk),
		.RCLKE(1),
		.RE(1),
		.WADDR(0),
		.WCLKN(0),
		.WCLKE(0),
		.WDATA(0),
		.WE(0)
		//.MASK(0) 
);

	SB_RAM512x8NRNW ram1(
		.RDATA(data_out_x[1][7:0]),
		.RADDR(addr_rd[8:0]),
		.RCLKN(clk),
		.RCLKE(1),
		.RE(1),
		.WADDR(0),
		.WCLKN(0),
		.WCLKE(0),
		.WDATA(0),
		.WE(0)
		//.MASK(0) 
);
	

endmodule
