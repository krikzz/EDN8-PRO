



module map_hub(
	input  MapIn mai,
	output MapOut mao
);

	
	
	
endmodule
