
module map_034(

	input  MapIn  mai,
	output MapOut mao
);
//************************************************************* base header
	CpuBus cpu;
	PpuBus ppu;
	SysCfg cfg;
	SSTBus sst;
	assign cpu = mai.cpu;
	assign ppu = mai.ppu;
	assign cfg = mai.cfg;
	assign sst = mai.sst;
	
	MemCtrl prg;
	MemCtrl chr;
	MemCtrl srm;
	assign mao.prg = prg;
	assign mao.chr = chr;
	assign mao.srm = srm;

	assign prg.dati			= cpu.data;
	assign chr.dati			= ppu.data;
	assign srm.dati			= cpu.data;
	
	wire int_cpu_oe;
	wire int_ppu_oe;
	wire [7:0]int_cpu_data;
	wire [7:0]int_ppu_data;
	
	assign mao.map_cpu_oe	= int_cpu_oe | (srm.ce & srm.oe) | (prg.ce & prg.oe);
	assign mao.map_cpu_do	= int_cpu_oe ? int_cpu_data : srm.ce ? mai.srm_do : mai.prg_do;
	
	assign mao.map_ppu_oe	= int_ppu_oe | (chr.ce & chr.oe);
	assign mao.map_ppu_do	= int_ppu_oe ? int_ppu_data : mai.chr_do;
//************************************************************* configuration
	assign mao.prg_mask_off = 0;
	assign mao.chr_mask_off = 0;
	assign mao.srm_mask_off = 0;
	assign mao.mir_4sc		= 0;//enable support for 4-screen mirroring. for activation should be enabled in cfg.mir_4 also
	assign mao.bus_cf 		= 0;//bus conflicts
//************************************************************* save state regs read
	assign mao.sst_di[7:0] =
	sst.addr[7:0] == 0 ? prg_reg : 
	sst.addr[7:0] == 1 ? chr0 : 
	sst.addr[7:0] == 2 ? chr1 : 
	sst.addr[7:0] == 127 ? cfg.map_idx : 8'hff;
//************************************************************* mapper-controlled pins
	assign srm.ce				= {cpu.addr[15:13], 13'd0} == 16'h6000;
	assign srm.oe				= cpu.rw;
	assign srm.we				= !cpu.rw;
	assign srm.addr[12:0]	= cpu.addr[12:0];
	
	assign prg.ce				= cpu.addr[15];
	assign prg.oe 				= cpu.rw;
	assign prg.we				= 0;
	assign prg.addr[14:0]	= cpu.addr[14:0];
	assign prg.addr[18:15] 	= !cpu.addr[15] ? 0 : prg_reg[3:0];
	
	assign chr.ce 				= mao.ciram_ce;
	assign chr.oe 				= !ppu.oe;
	assign chr.we 				= cfg.chr_ram ? !ppu.we & mao.ciram_ce : 0;
	assign chr.addr[11:0]	= ppu.addr[11:0];
	assign chr.addr[12] 		= cfg.chr_ram ? ppu.addr[12] : chr_reg[0];
	assign chr.addr[16:13] 	= chr_reg[4:1];

	
	//A10-Vmir, A11-Hmir
	assign mao.ciram_a10 	= cfg.mir_v ? ppu.addr[10] : ppu.addr[11];
	assign mao.ciram_ce 		= !ppu.addr[13];
	
	assign mao.irq				= 0;
//************************************************************* mapper implementation
	
	reg [3:0]prg_reg;
	reg [4:0]chr0;
	reg [4:0]chr1;
	
	wire [4:0]chr_reg = !ppu.addr[12] ? chr0[4:0] : chr1[4:0];
	
	always @(negedge cpu.m2)
	if(sst.act)
	begin
		if(sst.we_reg & sst.addr[7:0] == 0)prg_reg 	<= sst.dato[1:0];
		if(sst.we_reg & sst.addr[7:0] == 1)chr0 		<= sst.dato[1:0];
		if(sst.we_reg & sst.addr[7:0] == 2)chr1 		<= sst.dato[1:0];
	end
		else
	if(mai.map_rst)
	begin
		prg_reg <= 0;
	end
		else
	if(cfg.chr_ram == 1 & cpu.addr[15] == 1 & !cpu.rw)
	begin
		prg_reg[3:0] <= cpu.data[3:0];
	end
		else
	if(cfg.chr_ram == 0 & cpu.addr[15] == 0 & !cpu.rw)
	begin
		if(cpu.addr[14:0] == 15'h7FFD)prg_reg[3:0] 	<= cpu.data[3:0];
			else
		if(cpu.addr[14:0] == 15'h7FFE)chr0[4:0] 		<= cpu.data[4:0];
			else
		if(cpu.addr[14:0] == 15'h7FFF)chr1[4:0] 		<= cpu.data[4:0];
	end

	
endmodule
