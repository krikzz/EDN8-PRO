

	`define SST_ON	//remove save state
	`define GGC_ON	//remove cheats engine
	`define SND_ON	//remove expansion sound if any exists
