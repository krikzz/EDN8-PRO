module ym2413_exp_rom(a,d);

	input [7:0]		a;
	output reg [9:0]	d;
	
	always @* begin
		case (a[7:0])
			8'd0 : d = 10'd0;
			8'd1 : d = 10'd3;
			8'd2 : d = 10'd6;
			8'd3 : d = 10'd8;
			8'd4 : d = 10'd11;
			8'd5 : d = 10'd14;
			8'd6 : d = 10'd17;
			8'd7 : d = 10'd20;
			8'd8 : d = 10'd22;
			8'd9 : d = 10'd25;
			8'd10 : d = 10'd28;
			8'd11 : d = 10'd31;
			8'd12 : d = 10'd34;
			8'd13 : d = 10'd37;
			8'd14 : d = 10'd40;
			8'd15 : d = 10'd42;
			8'd16 : d = 10'd45;
			8'd17 : d = 10'd48;
			8'd18 : d = 10'd51;
			8'd19 : d = 10'd54;
			8'd20 : d = 10'd57;
			8'd21 : d = 10'd60;
			8'd22 : d = 10'd63;
			8'd23 : d = 10'd66;
			8'd24 : d = 10'd69;
			8'd25 : d = 10'd72;
			8'd26 : d = 10'd75;
			8'd27 : d = 10'd78;
			8'd28 : d = 10'd81;
			8'd29 : d = 10'd84;
			8'd30 : d = 10'd87;
			8'd31 : d = 10'd90;
			8'd32 : d = 10'd93;
			8'd33 : d = 10'd96;
			8'd34 : d = 10'd99;
			8'd35 : d = 10'd102;
			8'd36 : d = 10'd105;
			8'd37 : d = 10'd108;
			8'd38 : d = 10'd111;
			8'd39 : d = 10'd114;
			8'd40 : d = 10'd117;
			8'd41 : d = 10'd120;
			8'd42 : d = 10'd123;
			8'd43 : d = 10'd126;
			8'd44 : d = 10'd130;
			8'd45 : d = 10'd133;
			8'd46 : d = 10'd136;
			8'd47 : d = 10'd139;
			8'd48 : d = 10'd142;
			8'd49 : d = 10'd145;
			8'd50 : d = 10'd148;
			8'd51 : d = 10'd152;
			8'd52 : d = 10'd155;
			8'd53 : d = 10'd158;
			8'd54 : d = 10'd161;
			8'd55 : d = 10'd164;
			8'd56 : d = 10'd168;
			8'd57 : d = 10'd171;
			8'd58 : d = 10'd174;
			8'd59 : d = 10'd177;
			8'd60 : d = 10'd181;
			8'd61 : d = 10'd184;
			8'd62 : d = 10'd187;
			8'd63 : d = 10'd190;
			8'd64 : d = 10'd194;
			8'd65 : d = 10'd197;
			8'd66 : d = 10'd200;
			8'd67 : d = 10'd204;
			8'd68 : d = 10'd207;
			8'd69 : d = 10'd210;
			8'd70 : d = 10'd214;
			8'd71 : d = 10'd217;
			8'd72 : d = 10'd220;
			8'd73 : d = 10'd224;
			8'd74 : d = 10'd227;
			8'd75 : d = 10'd231;
			8'd76 : d = 10'd234;
			8'd77 : d = 10'd237;
			8'd78 : d = 10'd241;
			8'd79 : d = 10'd244;
			8'd80 : d = 10'd248;
			8'd81 : d = 10'd251;
			8'd82 : d = 10'd255;
			8'd83 : d = 10'd258;
			8'd84 : d = 10'd262;
			8'd85 : d = 10'd265;
			8'd86 : d = 10'd268;
			8'd87 : d = 10'd272;
			8'd88 : d = 10'd276;
			8'd89 : d = 10'd279;
			8'd90 : d = 10'd283;
			8'd91 : d = 10'd286;
			8'd92 : d = 10'd290;
			8'd93 : d = 10'd293;
			8'd94 : d = 10'd297;
			8'd95 : d = 10'd300;
			8'd96 : d = 10'd304;
			8'd97 : d = 10'd308;
			8'd98 : d = 10'd311;
			8'd99 : d = 10'd315;
			8'd100 : d = 10'd318;
			8'd101 : d = 10'd322;
			8'd102 : d = 10'd326;
			8'd103 : d = 10'd329;
			8'd104 : d = 10'd333;
			8'd105 : d = 10'd337;
			8'd106 : d = 10'd340;
			8'd107 : d = 10'd344;
			8'd108 : d = 10'd348;
			8'd109 : d = 10'd352;
			8'd110 : d = 10'd355;
			8'd111 : d = 10'd359;
			8'd112 : d = 10'd363;
			8'd113 : d = 10'd367;
			8'd114 : d = 10'd370;
			8'd115 : d = 10'd374;
			8'd116 : d = 10'd378;
			8'd117 : d = 10'd382;
			8'd118 : d = 10'd385;
			8'd119 : d = 10'd389;
			8'd120 : d = 10'd393;
			8'd121 : d = 10'd397;
			8'd122 : d = 10'd401;
			8'd123 : d = 10'd405;
			8'd124 : d = 10'd409;
			8'd125 : d = 10'd412;
			8'd126 : d = 10'd416;
			8'd127 : d = 10'd420;
			8'd128 : d = 10'd424;
			8'd129 : d = 10'd428;
			8'd130 : d = 10'd432;
			8'd131 : d = 10'd436;
			8'd132 : d = 10'd440;
			8'd133 : d = 10'd444;
			8'd134 : d = 10'd448;
			8'd135 : d = 10'd452;
			8'd136 : d = 10'd456;
			8'd137 : d = 10'd460;
			8'd138 : d = 10'd464;
			8'd139 : d = 10'd468;
			8'd140 : d = 10'd472;
			8'd141 : d = 10'd476;
			8'd142 : d = 10'd480;
			8'd143 : d = 10'd484;
			8'd144 : d = 10'd488;
			8'd145 : d = 10'd492;
			8'd146 : d = 10'd496;
			8'd147 : d = 10'd501;
			8'd148 : d = 10'd505;
			8'd149 : d = 10'd509;
			8'd150 : d = 10'd513;
			8'd151 : d = 10'd517;
			8'd152 : d = 10'd521;
			8'd153 : d = 10'd526;
			8'd154 : d = 10'd530;
			8'd155 : d = 10'd534;
			8'd156 : d = 10'd538;
			8'd157 : d = 10'd542;
			8'd158 : d = 10'd547;
			8'd159 : d = 10'd551;
			8'd160 : d = 10'd555;
			8'd161 : d = 10'd560;
			8'd162 : d = 10'd564;
			8'd163 : d = 10'd568;
			8'd164 : d = 10'd572;
			8'd165 : d = 10'd577;
			8'd166 : d = 10'd581;
			8'd167 : d = 10'd585;
			8'd168 : d = 10'd590;
			8'd169 : d = 10'd594;
			8'd170 : d = 10'd599;
			8'd171 : d = 10'd603;
			8'd172 : d = 10'd607;
			8'd173 : d = 10'd612;
			8'd174 : d = 10'd616;
			8'd175 : d = 10'd621;
			8'd176 : d = 10'd625;
			8'd177 : d = 10'd630;
			8'd178 : d = 10'd634;
			8'd179 : d = 10'd639;
			8'd180 : d = 10'd643;
			8'd181 : d = 10'd648;
			8'd182 : d = 10'd652;
			8'd183 : d = 10'd657;
			8'd184 : d = 10'd661;
			8'd185 : d = 10'd666;
			8'd186 : d = 10'd670;
			8'd187 : d = 10'd675;
			8'd188 : d = 10'd680;
			8'd189 : d = 10'd684;
			8'd190 : d = 10'd689;
			8'd191 : d = 10'd693;
			8'd192 : d = 10'd698;
			8'd193 : d = 10'd703;
			8'd194 : d = 10'd708;
			8'd195 : d = 10'd712;
			8'd196 : d = 10'd717;
			8'd197 : d = 10'd722;
			8'd198 : d = 10'd726;
			8'd199 : d = 10'd731;
			8'd200 : d = 10'd736;
			8'd201 : d = 10'd741;
			8'd202 : d = 10'd745;
			8'd203 : d = 10'd750;
			8'd204 : d = 10'd755;
			8'd205 : d = 10'd760;
			8'd206 : d = 10'd765;
			8'd207 : d = 10'd770;
			8'd208 : d = 10'd774;
			8'd209 : d = 10'd779;
			8'd210 : d = 10'd784;
			8'd211 : d = 10'd789;
			8'd212 : d = 10'd794;
			8'd213 : d = 10'd799;
			8'd214 : d = 10'd804;
			8'd215 : d = 10'd809;
			8'd216 : d = 10'd814;
			8'd217 : d = 10'd819;
			8'd218 : d = 10'd824;
			8'd219 : d = 10'd829;
			8'd220 : d = 10'd834;
			8'd221 : d = 10'd839;
			8'd222 : d = 10'd844;
			8'd223 : d = 10'd849;
			8'd224 : d = 10'd854;
			8'd225 : d = 10'd859;
			8'd226 : d = 10'd864;
			8'd227 : d = 10'd869;
			8'd228 : d = 10'd874;
			8'd229 : d = 10'd880;
			8'd230 : d = 10'd885;
			8'd231 : d = 10'd890;
			8'd232 : d = 10'd895;
			8'd233 : d = 10'd900;
			8'd234 : d = 10'd906;
			8'd235 : d = 10'd911;
			8'd236 : d = 10'd916;
			8'd237 : d = 10'd921;
			8'd238 : d = 10'd927;
			8'd239 : d = 10'd932;
			8'd240 : d = 10'd937;
			8'd241 : d = 10'd942;
			8'd242 : d = 10'd948;
			8'd243 : d = 10'd953;
			8'd244 : d = 10'd959;
			8'd245 : d = 10'd964;
			8'd246 : d = 10'd969;
			8'd247 : d = 10'd975;
			8'd248 : d = 10'd980;
			8'd249 : d = 10'd986;
			8'd250 : d = 10'd991;
			8'd251 : d = 10'd996;
			8'd252 : d = 10'd1002;
			8'd253 : d = 10'd1007;
			8'd254 : d = 10'd1013;
			8'd255 : d = 10'd1018;		
		endcase
	end
endmodule

module ym2413_logsin_rom(a,d);

	input [7:0]	a;
	output reg [11:0]	d;
	
	always @* begin
		case (a[7:0])	
			8'd0 : d = 12'd2137;
			8'd1 : d = 12'd1731;
			8'd2 : d = 12'd1543;
			8'd3 : d = 12'd1419;
			8'd4 : d = 12'd1326;
			8'd5 : d = 12'd1252;
			8'd6 : d = 12'd1190;
			8'd7 : d = 12'd1137;
			8'd8 : d = 12'd1091;
			8'd9 : d = 12'd1050;
			8'd10 : d = 12'd1013;
			8'd11 : d = 12'd979;
			8'd12 : d = 12'd949;
			8'd13 : d = 12'd920;
			8'd14 : d = 12'd894;
			8'd15 : d = 12'd869;
			8'd16 : d = 12'd846;
			8'd17 : d = 12'd825;
			8'd18 : d = 12'd804;
			8'd19 : d = 12'd785;
			8'd20 : d = 12'd767;
			8'd21 : d = 12'd749;
			8'd22 : d = 12'd732;
			8'd23 : d = 12'd717;
			8'd24 : d = 12'd701;
			8'd25 : d = 12'd687;
			8'd26 : d = 12'd672;
			8'd27 : d = 12'd659;
			8'd28 : d = 12'd646;
			8'd29 : d = 12'd633;
			8'd30 : d = 12'd621;
			8'd31 : d = 12'd609;
			8'd32 : d = 12'd598;
			8'd33 : d = 12'd587;
			8'd34 : d = 12'd576;
			8'd35 : d = 12'd566;
			8'd36 : d = 12'd556;
			8'd37 : d = 12'd546;
			8'd38 : d = 12'd536;
			8'd39 : d = 12'd527;
			8'd40 : d = 12'd518;
			8'd41 : d = 12'd509;
			8'd42 : d = 12'd501;
			8'd43 : d = 12'd492;
			8'd44 : d = 12'd484;
			8'd45 : d = 12'd476;
			8'd46 : d = 12'd468;
			8'd47 : d = 12'd461;
			8'd48 : d = 12'd453;
			8'd49 : d = 12'd446;
			8'd50 : d = 12'd439;
			8'd51 : d = 12'd432;
			8'd52 : d = 12'd425;
			8'd53 : d = 12'd418;
			8'd54 : d = 12'd411;
			8'd55 : d = 12'd405;
			8'd56 : d = 12'd399;
			8'd57 : d = 12'd392;
			8'd58 : d = 12'd386;
			8'd59 : d = 12'd380;
			8'd60 : d = 12'd375;
			8'd61 : d = 12'd369;
			8'd62 : d = 12'd363;
			8'd63 : d = 12'd358;
			8'd64 : d = 12'd352;
			8'd65 : d = 12'd347;
			8'd66 : d = 12'd341;
			8'd67 : d = 12'd336;
			8'd68 : d = 12'd331;
			8'd69 : d = 12'd326;
			8'd70 : d = 12'd321;
			8'd71 : d = 12'd316;
			8'd72 : d = 12'd311;
			8'd73 : d = 12'd307;
			8'd74 : d = 12'd302;
			8'd75 : d = 12'd297;
			8'd76 : d = 12'd293;
			8'd77 : d = 12'd289;
			8'd78 : d = 12'd284;
			8'd79 : d = 12'd280;
			8'd80 : d = 12'd276;
			8'd81 : d = 12'd271;
			8'd82 : d = 12'd267;
			8'd83 : d = 12'd263;
			8'd84 : d = 12'd259;
			8'd85 : d = 12'd255;
			8'd86 : d = 12'd251;
			8'd87 : d = 12'd248;
			8'd88 : d = 12'd244;
			8'd89 : d = 12'd240;
			8'd90 : d = 12'd236;
			8'd91 : d = 12'd233;
			8'd92 : d = 12'd229;
			8'd93 : d = 12'd226;
			8'd94 : d = 12'd222;
			8'd95 : d = 12'd219;
			8'd96 : d = 12'd215;
			8'd97 : d = 12'd212;
			8'd98 : d = 12'd209;
			8'd99 : d = 12'd205;
			8'd100 : d = 12'd202;
			8'd101 : d = 12'd199;
			8'd102 : d = 12'd196;
			8'd103 : d = 12'd193;
			8'd104 : d = 12'd190;
			8'd105 : d = 12'd187;
			8'd106 : d = 12'd184;
			8'd107 : d = 12'd181;
			8'd108 : d = 12'd178;
			8'd109 : d = 12'd175;
			8'd110 : d = 12'd172;
			8'd111 : d = 12'd169;
			8'd112 : d = 12'd167;
			8'd113 : d = 12'd164;
			8'd114 : d = 12'd161;
			8'd115 : d = 12'd159;
			8'd116 : d = 12'd156;
			8'd117 : d = 12'd153;
			8'd118 : d = 12'd151;
			8'd119 : d = 12'd148;
			8'd120 : d = 12'd146;
			8'd121 : d = 12'd143;
			8'd122 : d = 12'd141;
			8'd123 : d = 12'd138;
			8'd124 : d = 12'd136;
			8'd125 : d = 12'd134;
			8'd126 : d = 12'd131;
			8'd127 : d = 12'd129;
			8'd128 : d = 12'd127;
			8'd129 : d = 12'd125;
			8'd130 : d = 12'd122;
			8'd131 : d = 12'd120;
			8'd132 : d = 12'd118;
			8'd133 : d = 12'd116;
			8'd134 : d = 12'd114;
			8'd135 : d = 12'd112;
			8'd136 : d = 12'd110;
			8'd137 : d = 12'd108;
			8'd138 : d = 12'd106;
			8'd139 : d = 12'd104;
			8'd140 : d = 12'd102;
			8'd141 : d = 12'd100;
			8'd142 : d = 12'd98;
			8'd143 : d = 12'd96;
			8'd144 : d = 12'd94;
			8'd145 : d = 12'd92;
			8'd146 : d = 12'd91;
			8'd147 : d = 12'd89;
			8'd148 : d = 12'd87;
			8'd149 : d = 12'd85;
			8'd150 : d = 12'd83;
			8'd151 : d = 12'd82;
			8'd152 : d = 12'd80;
			8'd153 : d = 12'd78;
			8'd154 : d = 12'd77;
			8'd155 : d = 12'd75;
			8'd156 : d = 12'd74;
			8'd157 : d = 12'd72;
			8'd158 : d = 12'd70;
			8'd159 : d = 12'd69;
			8'd160 : d = 12'd67;
			8'd161 : d = 12'd66;
			8'd162 : d = 12'd64;
			8'd163 : d = 12'd63;
			8'd164 : d = 12'd62;
			8'd165 : d = 12'd60;
			8'd166 : d = 12'd59;
			8'd167 : d = 12'd57;
			8'd168 : d = 12'd56;
			8'd169 : d = 12'd55;
			8'd170 : d = 12'd53;
			8'd171 : d = 12'd52;
			8'd172 : d = 12'd51;
			8'd173 : d = 12'd49;
			8'd174 : d = 12'd48;
			8'd175 : d = 12'd47;
			8'd176 : d = 12'd46;
			8'd177 : d = 12'd45;
			8'd178 : d = 12'd43;
			8'd179 : d = 12'd42;
			8'd180 : d = 12'd41;
			8'd181 : d = 12'd40;
			8'd182 : d = 12'd39;
			8'd183 : d = 12'd38;
			8'd184 : d = 12'd37;
			8'd185 : d = 12'd36;
			8'd186 : d = 12'd35;
			8'd187 : d = 12'd34;
			8'd188 : d = 12'd33;
			8'd189 : d = 12'd32;
			8'd190 : d = 12'd31;
			8'd191 : d = 12'd30;
			8'd192 : d = 12'd29;
			8'd193 : d = 12'd28;
			8'd194 : d = 12'd27;
			8'd195 : d = 12'd26;
			8'd196 : d = 12'd25;
			8'd197 : d = 12'd24;
			8'd198 : d = 12'd23;
			8'd199 : d = 12'd23;
			8'd200 : d = 12'd22;
			8'd201 : d = 12'd21;
			8'd202 : d = 12'd20;
			8'd203 : d = 12'd20;
			8'd204 : d = 12'd19;
			8'd205 : d = 12'd18;
			8'd206 : d = 12'd17;
			8'd207 : d = 12'd17;
			8'd208 : d = 12'd16;
			8'd209 : d = 12'd15;
			8'd210 : d = 12'd15;
			8'd211 : d = 12'd14;
			8'd212 : d = 12'd13;
			8'd213 : d = 12'd13;
			8'd214 : d = 12'd12;
			8'd215 : d = 12'd12;
			8'd216 : d = 12'd11;
			8'd217 : d = 12'd10;
			8'd218 : d = 12'd10;
			8'd219 : d = 12'd9;
			8'd220 : d = 12'd9;
			8'd221 : d = 12'd8;
			8'd222 : d = 12'd8;
			8'd223 : d = 12'd7;
			8'd224 : d = 12'd7;
			8'd225 : d = 12'd7;
			8'd226 : d = 12'd6;
			8'd227 : d = 12'd6;
			8'd228 : d = 12'd5;
			8'd229 : d = 12'd5;
			8'd230 : d = 12'd5;
			8'd231 : d = 12'd4;
			8'd232 : d = 12'd4;
			8'd233 : d = 12'd4;
			8'd234 : d = 12'd3;
			8'd235 : d = 12'd3;
			8'd236 : d = 12'd3;
			8'd237 : d = 12'd2;
			8'd238 : d = 12'd2;
			8'd239 : d = 12'd2;
			8'd240 : d = 12'd2;
			8'd241 : d = 12'd1;
			8'd242 : d = 12'd1;
			8'd243 : d = 12'd1;
			8'd244 : d = 12'd1;
			8'd245 : d = 12'd1;
			8'd246 : d = 12'd1;
			8'd247 : d = 12'd1;
			8'd248 : d = 12'd0;
			8'd249 : d = 12'd0;
			8'd250 : d = 12'd0;
			8'd251 : d = 12'd0;
			8'd252 : d = 12'd0;
			8'd253 : d = 12'd0;
			8'd254 : d = 12'd0;
			8'd255 : d = 12'd0;
		endcase
	end

endmodule
