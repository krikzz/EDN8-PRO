

	`define SS_OFF	 	//remove save state
	`define GG_OFF	//remove cheats engine
	`define SND_OFF  //remove expansion sound if any exists
