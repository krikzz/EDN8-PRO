

	`define SST_OFF	//save state
	`define GGC_OFF	//cheats engine
	`define SND_OFF	//expansion sound if any exists
